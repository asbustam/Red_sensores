LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux_8a1vhdl IS
	
	PORT(DIN1:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		  DIN2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	
		  SEL:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		  DOUT:OUT STD_LOGIC_vector(7 DOWNTO 0));
	end mux_8a1vhdl ;

ARCHITECTURE BEH123 OF mux_8a1vhdl IS
BEGIN
PROCESS(DIN1,DIN2,SEL)
BEGIN
CASE SEL IS
WHEN"000"=>DOUT<="00100100";
WHEN"001"=>DOUT<="00000001";
WHEN"010"=>DOUT<="00000011";
WHEN"011"=>DOUT<=DIN1;
WHEN"100"=>DOUT<=DIN2;
WHEN"101"=>DOUT<="00000000";
WHEN"110"=>DOUT<="00000000";
WHEN"111"=>DOUT<="00000000";
--WHEN OTHERS=>DOUT<='ZZZZZZZZ';
END CASE;
END PROCESS;
END BEH123;