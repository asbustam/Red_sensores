LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY mux8a1 IS
	
PORT( A:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		B:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		C:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		D:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		E:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		F:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		G:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		H:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	   SEL:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	   Q:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END mux8a1 ;

ARCHITECTURE sol OF muX8a1 IS
BEGIN
	PROCESS(SEL,A,B,C,D,E,F,G,H)
	BEGIN
	CASE SEL IS
		WHEN"000"=>Q<=A;
		WHEN"001"=>Q<=B;
		WHEN"010"=>Q<="000000" & C;
		WHEN"011"=>Q<="0000" & D;
		WHEN"100"=>Q<=E;
		WHEN"101"=>Q<=F;
		WHEN"110"=>Q<=G;
		WHEN"111"=>Q<=H;
		WHEN OTHERS=>Q<="--------";
	END CASE;
	END PROCESS;
END sol;